//design(4'adder)

module adder(A,B,sum)

input A,B;
output sum;

assign sum = A+B;

endmodule